module simple_or(f,x,y);
	input x,y;
	output f;
	assign f=x|y;

endmodule
